// High level structural description language

#[VERSION_MIN "1.0"]
#[VERSION_MAX "1.0"]
#[VERSION_RECOMMENDED "1.0"]

#[PROJECT_NAME "Language Scratchpad"]
#[PROJECT_AUTHOR "John Earnest"]
#[PROJECT_DATE "2013-01-01"]

namespace storage::volatile
{
    primitive "sr_latch_gated"(set : line, en : line, reset : line)(q : line, qn : line)
    {
        tube S1, R1;

        on(reset)
        {
            S1 = 0;
            R1 = 1;
        }

        and(S1, en, set);
        and(R1, en, reset);
        nor(out, S1, q);
        nor(q, R1, qn);
    }

    template <int N>
    primitive "r"(set : line<N>, en : line, reset : line)(dat : line<N>)
    {
        basic sr_latch_gated bits[N];

        on(reset)
        {
            syncfor(i, 0, N)
            {
                bits[i].reset = 1;
            }
        }

        on(en)
        {
            syncfor(i, 0, N)
            {
                bits[i].en = 1;
            }

            syncfor(i, 0, N)
            {
                bits[i].set = set[i];
            }
        }

        syncfor(i, 0, N)
        {
            dat[i] = bits[i].q;
        }
    }

    // lets define 512 types of registers for sizes 1-512 inclusive
    metafor(i, 1, 512)
    {
        @/// @brief {{i}}-bit register primitive
        typedef r<{{i}}> r{{i}};
    }

    /// @brief SRAM primitive N size of width B
    template <int N, int W>
    primitive "static_ram_generic"(datin : line<W>, addr : line{{statics.math.log2(N)}}, writable : line, enable : line, reset : line)(dat : line<N>) : constraints(N > 0 && W > 0 && statics.math.ispow2(N))
    {
        basic r<W> regs[N];

        on(reset)
        {
            syncfor(i, 0, N)
            {
                regs[i].reset = 1;
            }
        }

        on(enable)
        {
            regs[addr].en = 1;

            on(writable)
            {
                regs[addr].set = datin;
            }

            dat = regs[addr].dat;
        }
    }
}

export module "sram_32K_8"(dat_in:line8, addr:line15, writable:line, enable:line, reset:line)(dat:line8)
{
    static_ram_generic<32768, 8> sram;

    sram.datin = dat_in;
    sram.addr = addr;
    sram.writable = writable;
    sram.enable = enable;
    sram.reset = reset;
}
